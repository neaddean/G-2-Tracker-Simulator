----------------------------------------------------------------------------------
-- function.vhd : convert binary to C5 code
--
-- inputs:
--   a     pulse number 0,1,2,3,4
--   B     C5 control or data code (0-15)
--   cd    '1' for control, '0' for data
--   q     '1' for Q0 (all normal pulses)
-- output:
--   Yout  four bit value to shift out LSB first to make the pulse
--
-- N.B. this is 100% combinatorial logic!
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
--use IEEE.STD_LOGIC_1076.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

entity funcgen is
  port (cd   : in  std_logic;
        a    : in  std_logic_vector(2 downto 0);  -- counter mod
        B    : in  std_logic_vector(3 downto 0);  -- code selector
        q0   : in  std_logic;                     -- send Q0
        Yout : out std_logic_vector (3 downto 0));
end funcgen;

architecture Behavioral of funcgen is
  signal inputs  : std_logic_vector (7 downto 0);
  signal outputs : std_logic_vector (1 downto 0);
begin

  inputs <= a & B & cd;
  with inputs select
    outputs <=
    "00" when "000" & "0000" & "0",     --D0
    "10" when "001" & "0000" & "0",
    "10" when "010" & "0000" & "0",
    "10" when "011" & "0000" & "0",
    "11" when "100" & "0000" & "0",

    "00" when "000" & "0001" & "0",     --D1
    "10" when "001" & "0001" & "0",
    "10" when "010" & "0001" & "0",
    "11" when "011" & "0001" & "0",
    "10" when "100" & "0001" & "0",

    "00" when "000" & "0010" & "0",     --D2
    "10" when "001" & "0010" & "0",
    "11" when "010" & "0010" & "0",
    "10" when "011" & "0010" & "0",
    "10" when "100" & "0010" & "0",

    "00" when "000" & "0011" & "0",     --D3
    "10" when "001" & "0011" & "0",
    "11" when "010" & "0011" & "0",
    "00" when "011" & "0011" & "0",
    "11" when "100" & "0011" & "0",

    "00" when "000" & "0100" & "0",     --D4
    "11" when "001" & "0100" & "0",
    "10" when "010" & "0100" & "0",
    "10" when "011" & "0100" & "0",
    "10" when "100" & "0100" & "0",

    "00" when "000" & "0101" & "0",     --D5
    "11" when "001" & "0101" & "0",
    "10" when "010" & "0101" & "0",
    "00" when "011" & "0101" & "0",
    "11" when "100" & "0101" & "0",

    "00" when "000" & "0110" & "0",     --D6
    "11" when "001" & "0110" & "0",
    "00" when "010" & "0110" & "0",
    "10" when "011" & "0110" & "0",
    "11" when "100" & "0110" & "0",

    "00" when "000" & "0111" & "0",     --D7
    "11" when "001" & "0111" & "0",
    "00" when "010" & "0111" & "0",
    "11" when "011" & "0111" & "0",
    "10" when "100" & "0111" & "0",

    "11" when "000" & "1000" & "0",     --D8
    "10" when "001" & "1000" & "0",
    "10" when "010" & "1000" & "0",
    "10" when "011" & "1000" & "0",
    "00" when "100" & "1000" & "0",

    "11" when "000" & "1001" & "0",     --D9
    "10" when "001" & "1001" & "0",
    "10" when "010" & "1001" & "0",
    "00" when "011" & "1001" & "0",
    "10" when "100" & "1001" & "0",

    "11" when "000" & "1010" & "0",     --D10
    "10" when "001" & "1010" & "0",
    "00" when "010" & "1010" & "0",
    "10" when "011" & "1010" & "0",
    "10" when "100" & "1010" & "0",

    "11" when "000" & "1011" & "0",     --D11
    "10" when "001" & "1011" & "0",
    "00" when "010" & "1011" & "0",
    "11" when "011" & "1011" & "0",
    "00" when "100" & "1011" & "0",

    "11" when "000" & "1100" & "0",     --D12
    "00" when "001" & "1100" & "0",
    "10" when "010" & "1100" & "0",
    "10" when "011" & "1100" & "0",
    "10" when "100" & "1100" & "0",

    "11" when "000" & "1101" & "0",     --D13
    "00" when "001" & "1101" & "0",
    "10" when "010" & "1101" & "0",
    "11" when "011" & "1101" & "0",
    "00" when "100" & "1101" & "0",

    "11" when "000" & "1110" & "0",     --D14
    "00" when "001" & "1110" & "0",
    "11" when "010" & "1110" & "0",
    "10" when "011" & "1110" & "0",
    "00" when "100" & "1110" & "0",

    "11" when "000" & "1111" & "0",     --D15
    "00" when "001" & "1111" & "0",
    "11" when "010" & "1111" & "0",
    "00" when "011" & "1111" & "0",
    "10" when "100" & "1111" & "0",

---------------------------------------------------------------------------

    "00" when "000" & "0011" & "1",     --C3
    "10" when "001" & "0011" & "1",
    "11" when "010" & "0011" & "1",
    "11" when "011" & "0011" & "1",
    "00" when "100" & "0011" & "1",

    "00" when "000" & "0101" & "1",     --C5
    "11" when "001" & "0101" & "1",
    "00" when "010" & "0101" & "1",
    "11" when "011" & "0101" & "1",
    "10" when "100" & "0101" & "1",

    "00" when "000" & "0110" & "1",     --C6
    "11" when "001" & "0110" & "1",
    "11" when "010" & "0110" & "1",
    "10" when "011" & "0110" & "1",
    "00" when "100" & "0110" & "1",

    "00" when "000" & "0111" & "1",     --C7
    "11" when "001" & "0111" & "1",
    "11" when "010" & "0111" & "1",
    "00" when "011" & "0111" & "1",
    "10" when "100" & "0111" & "1",

    "11" when "000" & "1011" & "1",     --C11
    "10" when "001" & "1011" & "1",
    "00" when "010" & "1011" & "1",
    "00" when "011" & "1011" & "1",
    "11" when "100" & "1011" & "1",

    "11" when "000" & "1101" & "1",     --C13
    "00" when "001" & "1101" & "1",
    "10" when "010" & "1101" & "1",
    "00" when "011" & "1101" & "1",
    "11" when "100" & "1101" & "1",

    "11" when "000" & "1110" & "1",     --C14
    "00" when "001" & "1110" & "1",
    "00" when "010" & "1110" & "1",
    "10" when "011" & "1110" & "1",
    "11" when "100" & "1110" & "1",

    "11" when "000" & "1111" & "1",     --C15
    "00" when "001" & "1111" & "1",
    "00" when "010" & "1111" & "1",
    "11" when "011" & "1111" & "1",
    "10" when "100" & "1111" & "1",

-------------------------------------------------------------------------------

    "10" when "000" & "0000" & "1",     --Q0
    "10" when "001" & "0000" & "1",
    "10" when "010" & "0000" & "1",
    "10" when "011" & "0000" & "1",
    "10" when "100" & "0000" & "1",

    "10" when others;

  with q0 select
    Yout <=
    "1100"              when '1',
    '1' & outputs & '0' when others;

end Behavioral;
